module top_module( input in, output out );
    assign out = !in; //Logical NOT
    //assign out = ~in; //Bitwise NOT
endmodule
